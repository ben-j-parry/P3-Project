// instrmem.sv
// RISC-V program instructions Module
// Ver: 1.0
// Date: 22/11/22

//is this the same as program memory

//5 bit address
module instrmem #(parameter )


endmodule