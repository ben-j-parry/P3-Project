// instrmem.sv
// RISC-V  instruction memory Module
// Ver: 1.0
// Date: 25/11/22

//is this the same as program memory

//5 bit address
module instrmem #(parameter )


endmodule